module CTRLUNIT (
	
);
	
endmodule

/**
 * 
 */